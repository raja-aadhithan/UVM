package ram_pkg;
        import uvm_pkg::*;// import the uvm_pkg
        `include "uvm_macros.svh"// include the uvm_macros.svh
        `include "tb_defs.sv"// include the tb_defs.sv
        `include "write_xtn.sv"// include write_xtn.sv and short_xtn.sv
        `include "short_xtn.sv"
endpackage